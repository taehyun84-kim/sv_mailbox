`include "apb_sequence.sv"